module synth (

    	//////////// ADC //////////
	//output		          		ADC_CONVST,
	//output		          		ADC_DIN,
	//input 		          		ADC_DOUT,
	//output		          		ADC_SCLK,

	//////////// Audio //////////
	input 		          		AUD_ADCDAT,
	inout 		          		AUD_ADCLRCK,
	inout 		          		AUD_BCLK,
	output		          		AUD_DACDAT,
	inout 		          		AUD_DACLRCK,
	output		          		AUD_XCK,

	//////////// CLOCK //////////
	//input 		          		CLOCK2_50,
	//input 		          		CLOCK3_50,
	//input 		          		CLOCK4_50,
	input 		          		CLOCK_50,

	//////////// SDRAM //////////
	//output		    [12:0]		DRAM_ADDR,
	//output		     [1:0]		DRAM_BA,
	//output		          		DRAM_CAS_N,
	//output		          		DRAM_CKE,
	//output		          		DRAM_CLK,
	//output		          		DRAM_CS_N,
	//inout 		    [15:0]		DRAM_DQ,
	//output		          		DRAM_LDQM,
	//output		          		DRAM_RAS_N,
	//output		          		DRAM_UDQM,
	//output		          		DRAM_WE_N,

	//////////// I2C for Audio and Video-In //////////
	output		          		FPGA_I2C_SCLK,
	inout 		          		FPGA_I2C_SDAT,

	//////////// SEG7 //////////
	//output		     [6:0]		HEX0,
	//output		     [6:0]		HEX1,
	//output		     [6:0]		HEX2,
	//output		     [6:0]		HEX3,
	//output		     [6:0]		HEX4,
	//output		     [6:0]		HEX5,

	//////////// IR //////////
	//input 		          		IRDA_RXD,
	//output		          		IRDA_TXD,

	//////////// KEY //////////
	input 		     [3:0]		KEY,

	//////////// LED //////////
	output		reg     [9:0]		LEDR,

	//////////// PS2 //////////
	inout 		          		PS2_CLK,
	//inout 		          		PS2_CLK2,
	inout 		          		PS2_DAT,
	//inout 		          		PS2_DAT2,


	//////////// Video-In //////////
	//input 		          		TD_CLK27,
	//input 		     [7:0]		TD_DATA,
	//input 		          		TD_HS,
	//output		          		TD_RESET_N,
	//input 		          		TD_VS,

	//////////// VGA //////////
	//output		          		VGA_BLANK_N,
	//output		     [7:0]		VGA_B,
	//output		          		VGA_CLK,
	//output		     [7:0]		VGA_G,
	//output		          		VGA_HS,
	//output		     [7:0]		VGA_R,
	//output		          		VGA_SYNC_N,
	//output		          		VGA_VS,

	//////////// GPIO_0, GPIO_0 connect to GPIO Default //////////
	//inout 		    [35:0]		GPIO_0,

	//////////// GPIO_1, GPIO_1 connect to GPIO Default //////////
	//inout 		    [35:0]		GPIO_1

	//////////// SW //////////
	input 		     [9:0]		SW
	
	

	
	
);

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/


/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/
wire clk;
assign clk = CLOCK_50;
wire rst;
assign rst = KEY[0];
 
// Internal Wires
wire				audio_in_available;
wire		[31:0]	left_channel_audio_in;
wire		[31:0]	right_channel_audio_in;
reg				read_audio_in;

wire				audio_out_allowed;
reg		[31:0]	left_channel_audio_out;
reg		[31:0]	right_channel_audio_out;
wire				write_audio_out;



// Internal Registers


// State Machine Registers

/*****************************************************************************
 *                         Finite State Machine(s)                           *
 *****************************************************************************/


/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/
// Controlling which filter is applied
always@(*) begin
	// MicIn input or Tone Generator input
	if(SW[0] == 1'b1)
	begin
		right_channel_audio_out = left_channel_audio_in;
		left_channel_audio_out = right_channel_audio_in;
		read_audio_in = audio_in_available & readValid;
		LEDR = {10{1'b1}};
	end
	else
	begin
		right_channel_audio_out = tone;
		left_channel_audio_out = tone;
		read_audio_in = readValid;
		LEDR = {10{1'b0}};
	end
end

assign write_audio_out			= audio_in_available & audio_out_allowed;

/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/

Audio_Controller Audio_Controllers (
	// Inputs
	.CLOCK_50					(clk),
	.reset						(~rst),

	.clear_audio_in_memory		(),
	.read_audio_in				(read_audio_in),
	
	.clear_audio_out_memory		(),
	.left_channel_audio_out		(left_channel_audio_out),
	.right_channel_audio_out	(right_channel_audio_out),
	.write_audio_out			(write_audio_out),

	.AUD_ADCDAT					(AUD_ADCDAT),

	// Bidirectionals
	.AUD_BCLK					(AUD_BCLK),
	.AUD_ADCLRCK				(AUD_ADCLRCK),
	.AUD_DACLRCK				(AUD_DACLRCK),

	// Outputs
	.audio_in_available			(audio_in_available),
	.left_channel_audio_in		(left_channel_audio_in),
	.right_channel_audio_in		(right_channel_audio_in),

	.audio_out_allowed			(audio_out_allowed),

	.AUD_XCK					(AUD_XCK),
	.AUD_DACDAT					(AUD_DACDAT)
);

avconf #(.USE_MIC_INPUT(1)) avc (
	.FPGA_I2C_SCLK				(FPGA_I2C_SCLK),
	.FPGA_I2C_SDAT				(FPGA_I2C_SDAT),
	.CLOCK_50					(clk),
	.reset						(~rst)
);

wire readValid;

/*****************************************************************************
 *                             Logic Circuit                            *
 *****************************************************************************/

wire [31:0] tone;
// Frequency Generator - borrowed from someone elses code
toneGenerator t0(
	.selection(SW[9:6]), // selecting between different frequencies
	.clock(CLOCK_50),
	.Tone(tone),
	.readValid(readValid)
);

endmodule

/* Peter - This looks like a square wave generator */
module toneSynth(Counts, clock, Out, readValid);
	
	input clock;
	output signed [31:0] Out;
	input [18:0] Counts;
	output readValid;

	reg [18:0] Q;
	reg [11:0] enableCount;

	always@(posedge clock) 
	begin
		if(enableCount == 12'd0)
			enableCount <= 12'd1042;
		else
			enableCount <= enableCount - 1'b1;
	
		if(Q == 19'd0)
			Q <= Counts;
		else
			Q <= Q - 1'b1;	
	end

	assign Out = (Q > ((Counts + 1'd1) / 2'd2)? 32'd10000000: -32'd10000000);
	assign readValid = (enableCount == 12'd0)? 1'b1: 1'b0;

endmodule

/* selects different timing speeds */
module toneGenerator(
    input [3:0] selection,
    input clock,
    output signed [31:0] Tone,
    output readValid
);

    reg [3:0] Freq1;
    reg [3:0] Freq2;
    reg [18:0] counts;

    always @(*) begin
        case(selection [3:0])
            4'd0: begin // C2
                Freq1 = 4'd0; Freq2 = 4'd0;
                counts = 19'd764200; // lowest note
            end
            4'd1: begin // D2
                Freq1 = 4'd0; Freq2 = 4'd1;
                counts = 19'd680936;
            end
            4'd2: begin // E2
                Freq1 = 4'd0; Freq2 = 4'd2;
                counts = 19'd606920;
            end
            4'd3: begin // F2
                Freq1 = 4'd0; Freq2 = 4'd3;
                counts = 19'd572600;
            end
            4'd4: begin // G2
                Freq1 = 4'd0; Freq2 = 4'd4;
                counts = 19'd510208;
            end
            4'd5: begin // A2
                Freq1 = 4'd0; Freq2 = 4'd5;
                counts = 19'd454544;
            end
            4'd6: begin // B2
                Freq1 = 4'd0; Freq2 = 4'd6;
                counts = 19'd405488;
            end
            4'd7: begin // C3
                Freq1 = 4'd0; Freq2 = 4'd7;
                counts = 19'd382280;
            end
            4'd8: begin // D3
                Freq1 = 4'd0; Freq2 = 4'd8;
                counts = 19'd340360;
            end
            4'd9: begin // E3
                Freq1 = 4'd0; Freq2 = 4'd9;
                counts = 19'd303512;
            end
            4'd10: begin // F3
                Freq1 = 4'd1; Freq2 = 4'd0;
                counts = 19'd286256;
            end
            4'd11: begin // G3
                Freq1 = 4'd1; Freq2 = 4'd1;
                counts = 19'd255112;
            end
            4'd12: begin // A3
                Freq1 = 4'd1; Freq2 = 4'd2;
                counts = 19'd227272;
            end
            4'd13: begin // B3
                Freq1 = 4'd1; Freq2 = 4'd3;
                counts = 19'd201272;
            end
            4'd14: begin // C4
                Freq1 = 4'd1; Freq2 = 4'd4;
                counts = 19'd190872; // highest note
            end
            default: begin
                Freq1 = 4'd0; Freq2 = 4'd0;
                counts = 19'd764200; // default to C2
            end
        endcase
    end
	 




	 
	 
    // Instantiate the toneSynth module
    toneSynth t0(
        .Counts(counts),
        .clock(clock),
        .Out(Tone),
        .readValid(readValid)
    );


endmodule
